module traffic_light(clk,rst,pass,R,G,Y);
input clk,rst,pass;
output R,G,Y;

//write your code here

endmodule

